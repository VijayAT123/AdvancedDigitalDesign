//all combinational

module control_unit (

    
)
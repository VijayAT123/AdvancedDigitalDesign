module instruction_decode (input [31:0] inst, output inst_type) {

    
}